class mc_common;
	static bit flag;
endclass
