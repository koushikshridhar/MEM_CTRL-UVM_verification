package wb_pkg;
	`include "uvm_pkg.sv"//only comment for EDA sims
	import uvm_pkg::*;

	`include "wb_tx.sv"
	`include "wb_sqr.sv"
	`include "wb_cov.sv"
	`include "wb_drv.sv"
	`include "wb_mon.sv"
	`include "wb_agent.sv"
endpackage
