`include "uvm_pkg.sv"//only comment for EDA sims
import uvm_pkg::*;
