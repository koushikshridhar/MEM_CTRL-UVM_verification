import wb_pkg::*;
import mc_mem_pkg::*;
