// ----------------------------------------------------
//UVM sqr: wb_sqr
//----------------------------------------------------
typedef uvm_sequencer#(wb_tx) wb_sqr;